library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

ENTITY TestProject is
port(
	CLK 			: in std_logic;
	OUT_VECTOR 	: out std_logic_vector(6 downto 0)
);
end entity TestProject;

architecture arch of TestProject is
begin


end architecture arch;